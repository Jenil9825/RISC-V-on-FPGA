module Add_ALU_tb();

reg [31:0] PC_out, imm_gen;
wire [31:0] add_alu_out;

initial begin

end
endmodule